library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Donut is
	port (
		clock, reset, run : in std_logic;
		data_in : in std_logic_vector(7 downto 0);
		data_in2 : in std_logic_vector(7 downto 0);
		reports : out std_logic_vector(2-1 downto 0)
	);
end Donut;

architecture Structure of Donut is
	--------------------------
	-- Component Declarations
	--------------------------
	COMPONENT ste_sim_2x
		PORT
		(
			bitvector	:	in std_logic_vector(255 downto 0);
			bitvector2	:	in std_logic_vector(255 downto 0);
			char_in		:	in std_logic_vector(7 downto 0);
			char_in2		:	in std_logic_vector(7 downto 0);
			clock, reset, run		:	in std_logic;
			Enable	:	in std_logic;
			match		:	out std_logic
		);
	END COMPONENT;

	COMPONENT Counter
		GENERIC	(target : INTEGER := 8;
			at_target : INTEGER := 0);
		PORT	(clock : IN std_logic;
			Enable, Reset, run : IN std_logic;
--			q : OUT std_logic_vector(11 DOWNTO 0);
			match : OUT std_logic);
	END COMPONENT;
	--------------------------
	-- Signal Declarations
	--------------------------
	--- STEs
	signal bitvector1MERGED2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector1MERGED2_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable1MERGED2 : std_logic := '1';
	signal match1MERGED2 : std_logic := '0';
	
	signal bitvector2MERGED3 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector2MERGED3_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable2MERGED3 : std_logic := '0';
	signal match2MERGED3 : std_logic := '0';
	
	signal bitvector2MERGED6 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector2MERGED6_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable2MERGED6 : std_logic := '0';
	signal match2MERGED6 : std_logic := '0';
	
	signal bitvector3MERGED4 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector3MERGED4_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable3MERGED4 : std_logic := '0';
	signal match3MERGED4 : std_logic := '0';
	
	signal bitvector4MERGED5 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector4MERGED5_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable4MERGED5 : std_logic := '0';
	signal match4MERGED5 : std_logic := '0';
	
	signal bitvector5MERGEDreport_2x5 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector5MERGEDreport_2x5_2 : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal Enable5MERGEDreport_2x5 : std_logic := '0';
	signal match5MERGEDreport_2x5 : std_logic := '0';
	
	signal bitvector6MERGED7 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector6MERGED7_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable6MERGED7 : std_logic := '0';
	signal match6MERGED7 : std_logic := '0';
	
	signal bitvector7MERGED8 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector7MERGED8_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable7MERGED8 : std_logic := '0';
	signal match7MERGED8 : std_logic := '0';
	
	signal bitvector8MERGED3 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal bitvector8MERGED3_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	signal Enable8MERGED3 : std_logic := '0';
	signal match8MERGED3 : std_logic := '0';
	
	signal bitvectorstart_2x1MERGED1 : std_logic_vector(255 downto 0) := "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111";
	signal bitvectorstart_2x1MERGED1_2 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000";
	signal Enablestart_2x1MERGED1 : std_logic := '1';
	signal matchstart_2x1MERGED1 : std_logic := '0';
	
	--- ORs
	
	--- ANDs
	
	--- Counters


begin
	--- STEs
	-- 1MERGED2
	ste1MERGED2 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector1MERGED2,
			bitvector2=>bitvector1MERGED2_2,
			Enable=>Enable1MERGED2,
			match=>match1MERGED2,
			run=>run);

	-- 2MERGED3
	ste2MERGED3 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector2MERGED3,
			bitvector2=>bitvector2MERGED3_2,
			Enable=>Enable2MERGED3,
			match=>match2MERGED3,
			run=>run);

	Enable2MERGED3 <= matchstart_2x1MERGED1;
	-- 2MERGED6
	ste2MERGED6 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector2MERGED6,
			bitvector2=>bitvector2MERGED6_2,
			Enable=>Enable2MERGED6,
			match=>match2MERGED6,
			run=>run);

	Enable2MERGED6 <= matchstart_2x1MERGED1;
	-- 3MERGED4
	ste3MERGED4 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector3MERGED4,
			bitvector2=>bitvector3MERGED4_2,
			Enable=>Enable3MERGED4,
			match=>match3MERGED4,
			run=>run);

	Enable3MERGED4 <= match1MERGED2 OR match7MERGED8;
	-- 4MERGED5
	ste4MERGED5 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector4MERGED5,
			bitvector2=>bitvector4MERGED5_2,
			Enable=>Enable4MERGED5,
			match=>match4MERGED5,
			run=>run);

	reports(0) <= match4MERGED5;
	Enable4MERGED5 <= match8MERGED3 OR match2MERGED3;
	-- 5MERGEDreport_2x5
	ste5MERGEDreport_2x5 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector5MERGEDreport_2x5,
			bitvector2=>bitvector5MERGEDreport_2x5_2,
			Enable=>Enable5MERGEDreport_2x5,
			match=>match5MERGEDreport_2x5,
			run=>run);

	reports(1) <= match5MERGEDreport_2x5;
	Enable5MERGEDreport_2x5 <= match3MERGED4;
	-- 6MERGED7
	ste6MERGED7 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector6MERGED7,
			bitvector2=>bitvector6MERGED7_2,
			Enable=>Enable6MERGED7,
			match=>match6MERGED7,
			run=>run);

	Enable6MERGED7 <= match1MERGED2;
	-- 7MERGED8
	ste7MERGED8 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector7MERGED8,
			bitvector2=>bitvector7MERGED8_2,
			Enable=>Enable7MERGED8,
			match=>match7MERGED8,
			run=>run);

	Enable7MERGED8 <= match2MERGED6;
	-- 8MERGED3
	ste8MERGED3 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvector8MERGED3,
			bitvector2=>bitvector8MERGED3_2,
			Enable=>Enable8MERGED3,
			match=>match8MERGED3,
			run=>run);

	Enable8MERGED3 <= match6MERGED7;
	-- start_2x1MERGED1
	stestart_2x1MERGED1 : ste_sim_2x
	port map(char_in=>data_in,
			char_in2=>data_in2,
			clock=>clock,
			reset=>reset,
			bitvector=>bitvectorstart_2x1MERGED1,
			bitvector2=>bitvectorstart_2x1MERGED1_2,
			Enable=>Enablestart_2x1MERGED1,
			match=>matchstart_2x1MERGED1,
			run=>run);

	

	reset_n <= not reset;
	
	--- ORs
	
	--- ANDs
	--- Counters
end Structure;